module structs

pub struct SystemInstruction {
pub:
	parts []Part @[json: parts]
}
