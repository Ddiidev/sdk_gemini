module structs

pub enum Roles {
	user
	model
}
