module structs

pub struct SystemInstruction {
pub mut:
	parts []Part @[json: parts]
}
