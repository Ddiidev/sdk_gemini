module structs

pub struct Part {
pub:
	text string @[json: text]
}
